library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

entity efinix_top is
    port (
        clock_120mhz : in std_logic;
        uart_rx      : in std_logic;
        uart_tx      : out std_logic
    );
end entity efinix_top;

architecture rtl of efinix_top is

    signal counter : integer range 0 to 2**16-1 := 0;

begin

    testi : process(clock_120mhz)
    begin
        if rising_edge(clock_120mhz) then
            if counter > 0 then
                counter <= counter - 1;
            else
                counter <= 1199;
                uart_tx <= uart_rx;
            end if;
        end if; --rising_edge
    end process testi;	

--------------------------------------------------
    -- u_hvhdl_example : entity work.hvhdl_example_interconnect
    -- port map(
    --     system_clock => clock_120mhz,
    --     hvhdl_example_interconnect_FPGA_in.communications_FPGA_in.uart_FPGA_in.uart_transreceiver_FPGA_in.uart_rx_fpga_in.uart_rx      => uart_rx,
    --     hvhdl_example_interconnect_FPGA_out.communications_FPGA_out.uart_FPGA_out.uart_transreceiver_FPGA_out.uart_tx_fpga_out.uart_tx => uart_tx);

end rtl;
