library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

entity chebyshev is
    port (
        clk : in std_logic	;
        data_to_be_filtered : integer;
        filter_output : integer
    );
end entity chebyshev;

architecture rtl of chebyshev is


begin


end rtl;
